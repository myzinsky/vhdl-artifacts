library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity i2c_picture is
    PORT(
        addr       : in  unsigned(10 downto 0);
        output     : out std_logic_vector(7 downto 0)
    );
end i2c_picture;

Architecture behavior of i2c_picture is

    type pixel is array (0 to 1023) of std_logic_vector(7 downto 0);
    signal picture : pixel := (
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00100000",
        "00100000",
        "00100000",
        "00100000",
        "00100000",
        "00100010",
        "00000010",
        "01000010",
        "01000010",
        "01000010",
        "01000000",
        "01000000",
        "00000000",
        "10000000",
        "10000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01100000",
        "00100000",
        "00110000",
        "00010000",
        "00010000",
        "00011000",
        "00001000",
        "10001000",
        "10001000",
        "10001100",
        "10000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "11000100",
        "10000100",
        "10000100",
        "10001100",
        "10001000",
        "10001000",
        "00001000",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "11000000",
        "01100000",
        "00110000",
        "00011000",
        "00001100",
        "10000100",
        "11000010",
        "11000010",
        "01100000",
        "00110000",
        "00011000",
        "00011000",
        "00001100",
        "10000100",
        "11000110",
        "11000010",
        "01100011",
        "00100011",
        "00110001",
        "00110001",
        "00010001",
        "00010000",
        "00011000",
        "10011000",
        "10011000",
        "10001000",
        "10001000",
        "10001000",
        "10001000",
        "10001000",
        "10001000",
        "10011000",
        "00011000",
        "00011000",
        "00010001",
        "00010001",
        "00110001",
        "00100001",
        "01100001",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000110",
        "00000011",
        "11000000",
        "01110000",
        "00111000",
        "00001100",
        "00000110",
        "10000011",
        "11100001",
        "00110000",
        "00011000",
        "00001100",
        "10000110",
        "11000011",
        "11100001",
        "01110001",
        "00111000",
        "00011000",
        "10011100",
        "10001100",
        "11000110",
        "11100110",
        "11100011",
        "01100011",
        "01110011",
        "00110011",
        "00110001",
        "00110001",
        "00110001",
        "00110001",
        "00110001",
        "00110001",
        "00110001",
        "00110001",
        "01110011",
        "01110011",
        "01100011",
        "11100010",
        "11000000",
        "11000000",
        "10000000",
        "00011000",
        "00011000",
        "00110000",
        "01110000",
        "11100000",
        "11000000",
        "10000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00001100",
        "00000111",
        "00000001",
        "11000000",
        "11110000",
        "00111100",
        "00001111",
        "00000011",
        "11100001",
        "11110000",
        "01111100",
        "00011110",
        "10001111",
        "11000111",
        "11110011",
        "01110001",
        "00111000",
        "00011100",
        "10001110",
        "11001110",
        "11100110",
        "11100111",
        "11100111",
        "01110111",
        "01110111",
        "01110111",
        "01100111",
        "11100111",
        "11100111",
        "11001110",
        "11001110",
        "10011100",
        "00011100",
        "01111000",
        "11110001",
        "11100011",
        "11000111",
        "00001110",
        "00011100",
        "01111000",
        "11110000",
        "11000011",
        "00000111",
        "00011110",
        "00111100",
        "00110000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011110",
        "00011111",
        "00000001",
        "00000000",
        "00010000",
        "00111111",
        "00011111",
        "00000001",
        "00000000",
        "00000100",
        "00000111",
        "00000111",
        "00000001",
        "00000000",
        "00001110",
        "00001111",
        "00001111",
        "00000011",
        "11111001",
        "11111100",
        "11111110",
        "00001110",
        "00001110",
        "00001110",
        "00011110",
        "11111100",
        "11111100",
        "11110001",
        "00000011",
        "00001111",
        "11111111",
        "11111100",
        "01000000",
        "00000011",
        "11111111",
        "11111111",
        "11111000",
        "00000000",
        "00000011",
        "11111111",
        "11111110",
        "00000000",
        "00000000",
        "00000000",
        "01111111",
        "00000100",
        "00000100",
        "00000100",
        "01111111",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00111000",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00101000",
        "00000000",
        "01111111",
        "00001000",
        "00000100",
        "00000100",
        "01111000",
        "00000000",
        "01001000",
        "01010100",
        "01010100",
        "01010100",
        "00100100",
        "00000000",
        "00111000",
        "01000100",
        "01000100",
        "01000100",
        "00101000",
        "00000000",
        "01111111",
        "00001000",
        "00000100",
        "00000100",
        "01111000",
        "00000000",
        "00111100",
        "01000000",
        "01000000",
        "01000000",
        "01111100",
        "00000000",
        "00111111",
        "01000000",
        "00000000",
        "00111000",
        "01010100",
        "01010100",
        "01010100",
        "01011000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00110000",
        "01110001",
        "01110011",
        "11100111",
        "11100111",
        "11100111",
        "11100111",
        "11100111",
        "11110111",
        "01110011",
        "01111001",
        "00111100",
        "00011111",
        "10001111",
        "11000011",
        "11110000",
        "01111100",
        "00111111",
        "00001111",
        "10000001",
        "11100000",
        "11111100",
        "00111111",
        "00001111",
        "00000000",
        "00000000",
        "00000000",
        "11000000",
        "00000000",
        "00000000",
        "10000000",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "11000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "10000000",
        "11000000",
        "10000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00001110",
        "00001110",
        "00001110",
        "00000111",
        "00000111",
        "00000011",
        "00000001",
        "00011000",
        "00011100",
        "00011110",
        "00001111",
        "11000111",
        "11100001",
        "01110000",
        "00111000",
        "00011110",
        "00000110",
        "00000000",
        "00000000",
        "00011111",
        "00000001",
        "00000001",
        "00000010",
        "00011100",
        "00000000",
        "00001000",
        "00010101",
        "00010101",
        "00010101",
        "00011110",
        "00000000",
        "00011111",
        "00000000",
        "00010010",
        "00010101",
        "00010101",
        "00010101",
        "00001001",
        "00000000",
        "00001110",
        "00010101",
        "00010101",
        "00010101",
        "00010110",
        "00000000",
        "00011111",
        "00000010",
        "00000001",
        "00000001",
        "00000010",
        "00000000",
        "00010010",
        "00010101",
        "00010101",
        "00010101",
        "00001001",
        "00000000",
        "00001111",
        "00010000",
        "00000000",
        "00001000",
        "00010101",
        "00010101",
        "00010101",
        "00011110",
        "00000000",
        "00001111",
        "00010000",
        "00010000",
        "00010000",
        "00011111",
        "00000000",
        "00000000",
        "00001111",
        "00010000",
        "00000000",
        "00001110",
        "00010101",
        "00010101",
        "00010101",
        "00010110",
        "00000000",
        "00011111",
        "00000010",
        "00000001",
        "00000001",
        "00000010",
        "00000000",
        "00011111",
        "00000001",
        "00000001",
        "00000001",
        "00011110",
        "00000000",
        "00000000"
    );  

begin

    output <= picture(to_integer(addr));

end behavior;
